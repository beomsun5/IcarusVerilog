module f_not(A, Q);
  // Input variable A
  input A;
  // Output variable Q
  output Q;
  assign Q = ~A;
endmodule